interface tx_intf(input WBCLK);
  logic        STX_PAD_O ;    // serial Transmitter output signal
  logic        BAUD_O;
endinterface: tx_intf
