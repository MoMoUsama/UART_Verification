package uart_agent_pkg;

  import uvm_pkg::*;
  import Env_Config_pkg::*;
  `include "uvm_macros.svh"

  `include "uart_seq_item.svh"
  `include "uart_driver.svh"
  `include "uart_monitor.svh"
  `include "uart_sequencer.svh"
  `include "uart_agent.svh"
  
endpackage : uart_agent_pkg
