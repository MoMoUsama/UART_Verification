interface rx_intf(input WBCLK);
  logic        SRX_PAD_I;    // serial Reciever input signal
endinterface: rx_intf