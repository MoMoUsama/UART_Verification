interface irq_intf;
  logic        INT_O ;    // Interrupt output signal
  
endinterface: irq_intf