package Env_Config_pkg;

  import uvm_pkg::*;
  `include "uvm_macros.svh"

  `include "ENV_Config.svh"
  
endpackage : Env_Config_pkg
